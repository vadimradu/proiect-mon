--driver pentru afisajul cu sapte segmente
